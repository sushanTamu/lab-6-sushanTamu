///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// Created by  : Prof. Quinn and Saumil Gogri
///////////////////////////////////////////////////////////////////////////


package htax_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "htax_packet_c.sv"
	`include "htax_sequencer_c.sv"
	`include "htax_tx_driver_c.svp"
	`include "htax_tx_agent_c.sv"
	`include "htax_seqs.sv"

endpackage
